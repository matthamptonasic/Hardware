/*
###############################################################################
#   Licensing information found at: 
#     https://github.com/hammy025/Hardware/
#   In file LICENSING.md
###############################################################################
#
#   File          :   dut.svh 
#   Creator       :   Matt Hampton (hammy025@gmail.com)
#   Owner         :   Matt Hampton (hammy025@gmail.com)
#   Creation Date :   04/05/16
#   Description   :   
#
###############################################################################
*/
`ifndef FIFO_FF_DUT_WIDTH
  `define FIFO_FF_DUT_WIDTH 32
`endif

`ifndef FIFO_FF_DUT_DEPTH
  `define FIFO_FF_DUT_DEPTH 16
`endif

