/*
###############################################################################
#   Licensing information found at: 
#     https://github.com/matthamptonasic/Hardware/
#   In file LICENSING.md
###############################################################################
#
#   File          :   dut.svh 
#   Creator       :   Matt Hampton (matthamptonasic@gmail.com)
#   Owner         :   Matt Hampton (matthamptonasic@gmail.com)
#   Creation Date :   04/05/16
#   Description   :   
#
###############################################################################
*/
`ifndef FIFO_FF_DUT_WIDTH
  `define FIFO_FF_DUT_WIDTH 32
`endif

`ifndef FIFO_FF_DUT_DEPTH
  `define FIFO_FF_DUT_DEPTH 16
`endif

